// nios_system.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                                            //                                       clk.clk
		input  wire        clk_0_clk,                                          //                                     clk_0.clk
		output wire [12:0] new_sdram_controller_0_wire_addr,                   //               new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,                     //                                          .ba
		output wire        new_sdram_controller_0_wire_cas_n,                  //                                          .cas_n
		output wire        new_sdram_controller_0_wire_cke,                    //                                          .cke
		output wire        new_sdram_controller_0_wire_cs_n,                   //                                          .cs_n
		inout  wire [31:0] new_sdram_controller_0_wire_dq,                     //                                          .dq
		output wire [3:0]  new_sdram_controller_0_wire_dqm,                    //                                          .dqm
		output wire        new_sdram_controller_0_wire_ras_n,                  //                                          .ras_n
		output wire        new_sdram_controller_0_wire_we_n,                   //                                          .we_n
		input  wire        reset_reset_n,                                      //                                     reset.reset_n
		input  wire        reset_0_reset_n,                                    //                                   reset_0.reset_n
		inout  wire [15:0] sram_0_external_interface_DQ,                       //                 sram_0_external_interface.DQ
		output wire [19:0] sram_0_external_interface_ADDR,                     //                                          .ADDR
		output wire        sram_0_external_interface_LB_N,                     //                                          .LB_N
		output wire        sram_0_external_interface_UB_N,                     //                                          .UB_N
		output wire        sram_0_external_interface_CE_N,                     //                                          .CE_N
		output wire        sram_0_external_interface_OE_N,                     //                                          .OE_N
		output wire        sram_0_external_interface_WE_N,                     //                                          .WE_N
		output wire [22:0] tristate_conduit_bridge_0_out_tcm_address_out,      //             tristate_conduit_bridge_0_out.tcm_address_out
		output wire [0:0]  tristate_conduit_bridge_0_out_tcm_read_n_out,       //                                          .tcm_read_n_out
		output wire [0:0]  tristate_conduit_bridge_0_out_tcm_write_n_out,      //                                          .tcm_write_n_out
		inout  wire [7:0]  tristate_conduit_bridge_0_out_tcm_data_out,         //                                          .tcm_data_out
		output wire [0:0]  tristate_conduit_bridge_0_out_tcm_chipselect_n_out, //                                          .tcm_chipselect_n_out
		output wire        video_vga_controller_0_external_interface_CLK,      // video_vga_controller_0_external_interface.CLK
		output wire        video_vga_controller_0_external_interface_HS,       //                                          .HS
		output wire        video_vga_controller_0_external_interface_VS,       //                                          .VS
		output wire        video_vga_controller_0_external_interface_BLANK,    //                                          .BLANK
		output wire        video_vga_controller_0_external_interface_SYNC,     //                                          .SYNC
		output wire [7:0]  video_vga_controller_0_external_interface_R,        //                                          .R
		output wire [7:0]  video_vga_controller_0_external_interface_G,        //                                          .G
		output wire [7:0]  video_vga_controller_0_external_interface_B         //                                          .B
	);

	wire         video_alpha_blender_0_avalon_blended_source_valid;                                        // video_alpha_blender_0:output_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] video_alpha_blender_0_avalon_blended_source_data;                                         // video_alpha_blender_0:output_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_alpha_blender_0_avalon_blended_source_ready;                                        // video_dual_clock_buffer_0:stream_in_ready -> video_alpha_blender_0:output_ready
	wire         video_alpha_blender_0_avalon_blended_source_startofpacket;                                // video_alpha_blender_0:output_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         video_alpha_blender_0_avalon_blended_source_endofpacket;                                  // video_alpha_blender_0:output_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_valid;                               // video_character_buffer_with_dma_0:stream_valid -> video_alpha_blender_0:foreground_valid
	wire  [39:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                // video_character_buffer_with_dma_0:stream_data -> video_alpha_blender_0:foreground_data
	wire         video_character_buffer_with_dma_0_avalon_char_source_ready;                               // video_alpha_blender_0:foreground_ready -> video_character_buffer_with_dma_0:stream_ready
	wire         video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                       // video_character_buffer_with_dma_0:stream_startofpacket -> video_alpha_blender_0:foreground_startofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                         // video_character_buffer_with_dma_0:stream_endofpacket -> video_alpha_blender_0:foreground_endofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                                  // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                                   // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                                  // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                          // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                            // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_valid;                                       // video_pixel_buffer_dma_0:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [15:0] video_pixel_buffer_dma_0_avalon_pixel_source_data;                                        // video_pixel_buffer_dma_0:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_ready;                                       // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma_0:stream_ready
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;                               // video_pixel_buffer_dma_0:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;                                 // video_pixel_buffer_dma_0:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                                            // video_rgb_resampler_0:stream_out_valid -> video_alpha_blender_0:background_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                             // video_rgb_resampler_0:stream_out_data -> video_alpha_blender_0:background_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                                            // video_alpha_blender_0:background_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                                    // video_rgb_resampler_0:stream_out_startofpacket -> video_alpha_blender_0:background_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                                      // video_rgb_resampler_0:stream_out_endofpacket -> video_alpha_blender_0:background_endofpacket
	wire         generic_tristate_controller_0_tcm_data_outen;                                             // generic_tristate_controller_0:tcm_data_outen -> tristate_conduit_bridge_0:tcs_tcm_data_outen
	wire         generic_tristate_controller_0_tcm_request;                                                // generic_tristate_controller_0:tcm_request -> tristate_conduit_bridge_0:request
	wire         generic_tristate_controller_0_tcm_write_n_out;                                            // generic_tristate_controller_0:tcm_write_n_out -> tristate_conduit_bridge_0:tcs_tcm_write_n_out
	wire         generic_tristate_controller_0_tcm_read_n_out;                                             // generic_tristate_controller_0:tcm_read_n_out -> tristate_conduit_bridge_0:tcs_tcm_read_n_out
	wire         generic_tristate_controller_0_tcm_grant;                                                  // tristate_conduit_bridge_0:grant -> generic_tristate_controller_0:tcm_grant
	wire         generic_tristate_controller_0_tcm_chipselect_n_out;                                       // generic_tristate_controller_0:tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_tcm_chipselect_n_out
	wire  [22:0] generic_tristate_controller_0_tcm_address_out;                                            // generic_tristate_controller_0:tcm_address_out -> tristate_conduit_bridge_0:tcs_tcm_address_out
	wire   [7:0] generic_tristate_controller_0_tcm_data_out;                                               // generic_tristate_controller_0:tcm_data_out -> tristate_conduit_bridge_0:tcs_tcm_data_out
	wire   [7:0] generic_tristate_controller_0_tcm_data_in;                                                // tristate_conduit_bridge_0:tcs_tcm_data_in -> generic_tristate_controller_0:tcm_data_in
	wire  [31:0] nios2_qsys_0_custom_instruction_master_result;                                            // nios2_qsys_0_custom_instruction_master_translator:ci_slave_result -> nios2_qsys_0:E_ci_combo_result
	wire         nios2_qsys_0_custom_instruction_master_readra;                                            // nios2_qsys_0:E_ci_combo_readra -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_qsys_0_custom_instruction_master_a;                                                 // nios2_qsys_0:E_ci_combo_a -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_qsys_0_custom_instruction_master_b;                                                 // nios2_qsys_0:E_ci_combo_b -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_c;                                                 // nios2_qsys_0:E_ci_combo_c -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_c
	wire         nios2_qsys_0_custom_instruction_master_readrb;                                            // nios2_qsys_0:E_ci_combo_readrb -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_readrb
	wire         nios2_qsys_0_custom_instruction_master_estatus;                                           // nios2_qsys_0:E_ci_combo_estatus -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_ipending;                                          // nios2_qsys_0:E_ci_combo_ipending -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_ipending
	wire  [31:0] nios2_qsys_0_custom_instruction_master_datab;                                             // nios2_qsys_0:E_ci_combo_datab -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_qsys_0_custom_instruction_master_dataa;                                             // nios2_qsys_0:E_ci_combo_dataa -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_writerc;                                           // nios2_qsys_0:E_ci_combo_writerc -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_writerc
	wire   [7:0] nios2_qsys_0_custom_instruction_master_n;                                                 // nios2_qsys_0:E_ci_combo_n -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_result;                  // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readra;                  // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_readra -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_a;                       // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_a -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_b;                       // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_b -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readrb;                  // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_c;                       // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_c -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_estatus;                 // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_ipending;                // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_datab;                   // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_datab -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_dataa;                   // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_writerc;                 // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_n;                       // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_n -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_result;                   // nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readra;                   // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_a;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_b;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readrb;                   // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_c;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_estatus;                  // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_ipending;                 // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_datab;                    // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_dataa;                    // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_writerc;                  // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_n;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_result;           // floating_point_adder_0:O -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_datab;            // nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_master_datab -> floating_point_adder_0:B
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa;            // nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> floating_point_adder_0:A
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_result;                   // nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_result -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_result
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_readra;                   // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_readra -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_a;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_a -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_a
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_b;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_b -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_b
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_readrb;                   // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_readrb -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_c;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_c -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_c
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_estatus;                  // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_estatus -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_ipending;                 // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_ipending -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_ipending
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_datab;                    // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_datab -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_dataa;                    // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_dataa -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_writerc;                  // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_writerc -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_writerc
	wire   [7:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_n;                        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master1_n -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_slave_n
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_result;           // floating_point_multiplier_0:O -> nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_master_result
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_datab;            // nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_master_datab -> floating_point_multiplier_0:B
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_dataa;            // nios2_qsys_0_custom_instruction_master_comb_slave_translator1:ci_master_dataa -> floating_point_multiplier_0:A
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;                             // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma_0:master_waitrequest
	wire  [15:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;                                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma_0:master_readdata
	wire  [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;                                 // video_pixel_buffer_dma_0:master_address -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_address
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;                                    // video_pixel_buffer_dma_0:master_read -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_read
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;                           // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma_0:master_readdatavalid
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock;                                    // video_pixel_buffer_dma_0:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                        // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                                     // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                                                     // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [28:0] nios2_qsys_0_data_master_address;                                                         // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                      // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                                            // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                                                   // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                                                           // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                       // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                 // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                                              // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                                                  // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                                                     // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                                            // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_readdata;                                      // sram_0:readdata -> mm_interconnect_0:sram_0_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_0_avalon_sram_slave_address;                                       // mm_interconnect_0:sram_0_avalon_sram_slave_address -> sram_0:address
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_read;                                          // mm_interconnect_0:sram_0_avalon_sram_slave_read -> sram_0:read
	wire   [1:0] mm_interconnect_0_sram_0_avalon_sram_slave_byteenable;                                    // mm_interconnect_0:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid;                                 // sram_0:readdatavalid -> mm_interconnect_0:sram_0_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_0_avalon_sram_slave_write;                                         // mm_interconnect_0:sram_0_avalon_sram_slave_write -> sram_0:write
	wire  [15:0] mm_interconnect_0_sram_0_avalon_sram_slave_writedata;                                     // mm_interconnect_0:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata;    // video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest; // video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address;     // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read;        // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata;   // video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address;    // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	wire   [3:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write;      // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata;                 // video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address;                  // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read;                     // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	wire   [3:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable;               // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write;                    // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata;                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                                 // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                              // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_readdata;                           // performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	wire   [4:0] mm_interconnect_0_performance_counter_0_control_slave_address;                            // mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_0_performance_counter_0_control_slave_begintransfer;                      // mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_0_performance_counter_0_control_slave_write;                              // mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_writedata;                          // mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;                                // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest;                             // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess;                             // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;                                 // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;                                    // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;                              // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;                                   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;                               // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;                                   // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;                                     // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;                                  // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;                                      // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;                                         // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [3:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;                                   // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;                                // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;                                        // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;                                    // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                                  // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                                    // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                                     // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                                       // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                                   // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [7:0] mm_interconnect_0_generic_tristate_controller_0_uas_readdata;                             // generic_tristate_controller_0:uas_readdata -> mm_interconnect_0:generic_tristate_controller_0_uas_readdata
	wire         mm_interconnect_0_generic_tristate_controller_0_uas_waitrequest;                          // generic_tristate_controller_0:uas_waitrequest -> mm_interconnect_0:generic_tristate_controller_0_uas_waitrequest
	wire         mm_interconnect_0_generic_tristate_controller_0_uas_debugaccess;                          // mm_interconnect_0:generic_tristate_controller_0_uas_debugaccess -> generic_tristate_controller_0:uas_debugaccess
	wire  [22:0] mm_interconnect_0_generic_tristate_controller_0_uas_address;                              // mm_interconnect_0:generic_tristate_controller_0_uas_address -> generic_tristate_controller_0:uas_address
	wire         mm_interconnect_0_generic_tristate_controller_0_uas_read;                                 // mm_interconnect_0:generic_tristate_controller_0_uas_read -> generic_tristate_controller_0:uas_read
	wire   [0:0] mm_interconnect_0_generic_tristate_controller_0_uas_byteenable;                           // mm_interconnect_0:generic_tristate_controller_0_uas_byteenable -> generic_tristate_controller_0:uas_byteenable
	wire         mm_interconnect_0_generic_tristate_controller_0_uas_readdatavalid;                        // generic_tristate_controller_0:uas_readdatavalid -> mm_interconnect_0:generic_tristate_controller_0_uas_readdatavalid
	wire         mm_interconnect_0_generic_tristate_controller_0_uas_lock;                                 // mm_interconnect_0:generic_tristate_controller_0_uas_lock -> generic_tristate_controller_0:uas_lock
	wire         mm_interconnect_0_generic_tristate_controller_0_uas_write;                                // mm_interconnect_0:generic_tristate_controller_0_uas_write -> generic_tristate_controller_0:uas_write
	wire   [7:0] mm_interconnect_0_generic_tristate_controller_0_uas_writedata;                            // mm_interconnect_0:generic_tristate_controller_0_uas_writedata -> generic_tristate_controller_0:uas_writedata
	wire   [0:0] mm_interconnect_0_generic_tristate_controller_0_uas_burstcount;                           // mm_interconnect_0:generic_tristate_controller_0_uas_burstcount -> generic_tristate_controller_0:uas_burstcount
	wire         irq_mapper_receiver0_irq;                                                                 // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                 // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                   // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                                                           // rst_controller:reset_out -> [generic_tristate_controller_0:reset_reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_qsys_0:reset_n, performance_counter_0:reset_n, rst_translator:in_reset, sram_0:reset, timer_0:reset_n, tristate_conduit_bridge_0:reset, video_alpha_blender_0:reset, video_character_buffer_with_dma_0:reset, video_dual_clock_buffer_0:reset_stream_in, video_pixel_buffer_dma_0:reset, video_rgb_resampler_0:reset]
	wire         rst_controller_reset_out_reset_req;                                                       // rst_controller:reset_req -> [nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                               // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                                       // rst_controller_001:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]

	fp_adder floating_point_adder_0 (
		.A (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.B (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //                              .datab
		.O (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_result)  //                              .result
	);

	fp_multiplier floating_point_multiplier_0 (
		.A (nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.B (nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_datab),  //                              .datab
		.O (nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_result)  //                              .result
	);

	nios_system_generic_tristate_controller_0 #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) generic_tristate_controller_0 (
		.clk_clk              (clk_clk),                                                           //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                                    // reset.reset
		.uas_address          (mm_interconnect_0_generic_tristate_controller_0_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_generic_tristate_controller_0_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_generic_tristate_controller_0_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_generic_tristate_controller_0_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_generic_tristate_controller_0_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_generic_tristate_controller_0_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_generic_tristate_controller_0_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_generic_tristate_controller_0_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_generic_tristate_controller_0_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_generic_tristate_controller_0_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_generic_tristate_controller_0_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (generic_tristate_controller_0_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (generic_tristate_controller_0_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (generic_tristate_controller_0_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (generic_tristate_controller_0_tcm_request),                         //      .request
		.tcm_grant            (generic_tristate_controller_0_tcm_grant),                           //      .grant
		.tcm_address_out      (generic_tristate_controller_0_tcm_address_out),                     //      .address_out
		.tcm_data_out         (generic_tristate_controller_0_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (generic_tristate_controller_0_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (generic_tristate_controller_0_tcm_data_in)                          //      .data_in
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                                                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                           //      .export
	);

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_combo_result                     (nios2_qsys_0_custom_instruction_master_result),                // custom_instruction_master.result
		.E_ci_combo_a                          (nios2_qsys_0_custom_instruction_master_a),                     //                          .a
		.E_ci_combo_b                          (nios2_qsys_0_custom_instruction_master_b),                     //                          .b
		.E_ci_combo_c                          (nios2_qsys_0_custom_instruction_master_c),                     //                          .c
		.E_ci_combo_dataa                      (nios2_qsys_0_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_combo_datab                      (nios2_qsys_0_custom_instruction_master_datab),                 //                          .datab
		.E_ci_combo_estatus                    (nios2_qsys_0_custom_instruction_master_estatus),               //                          .estatus
		.E_ci_combo_ipending                   (nios2_qsys_0_custom_instruction_master_ipending),              //                          .ipending
		.E_ci_combo_n                          (nios2_qsys_0_custom_instruction_master_n),                     //                          .n
		.E_ci_combo_readra                     (nios2_qsys_0_custom_instruction_master_readra),                //                          .readra
		.E_ci_combo_readrb                     (nios2_qsys_0_custom_instruction_master_readrb),                //                          .readrb
		.E_ci_combo_writerc                    (nios2_qsys_0_custom_instruction_master_writerc)                //                          .writerc
	);

	nios_system_performance_counter_0 performance_counter_0 (
		.clk           (clk_clk),                                                             //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                     //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	nios_system_sram_0 sram_0 (
		.clk           (clk_clk),                                                  //                clk.clk
		.reset         (rst_controller_reset_out_reset),                           //              reset.reset
		.SRAM_DQ       (sram_0_external_interface_DQ),                             // external_interface.export
		.SRAM_ADDR     (sram_0_external_interface_ADDR),                           //                   .export
		.SRAM_LB_N     (sram_0_external_interface_LB_N),                           //                   .export
		.SRAM_UB_N     (sram_0_external_interface_UB_N),                           //                   .export
		.SRAM_CE_N     (sram_0_external_interface_CE_N),                           //                   .export
		.SRAM_OE_N     (sram_0_external_interface_OE_N),                           //                   .export
		.SRAM_WE_N     (sram_0_external_interface_WE_N),                           //                   .export
		.address       (mm_interconnect_0_sram_0_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_0_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_0_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	nios_system_tristate_conduit_bridge_0 tristate_conduit_bridge_0 (
		.clk                      (clk_clk),                                            //   clk.clk
		.reset                    (rst_controller_reset_out_reset),                     // reset.reset
		.request                  (generic_tristate_controller_0_tcm_request),          //   tcs.request
		.grant                    (generic_tristate_controller_0_tcm_grant),            //      .grant
		.tcs_tcm_address_out      (generic_tristate_controller_0_tcm_address_out),      //      .address_out
		.tcs_tcm_read_n_out       (generic_tristate_controller_0_tcm_read_n_out),       //      .read_n_out
		.tcs_tcm_write_n_out      (generic_tristate_controller_0_tcm_write_n_out),      //      .write_n_out
		.tcs_tcm_data_out         (generic_tristate_controller_0_tcm_data_out),         //      .data_out
		.tcs_tcm_data_outen       (generic_tristate_controller_0_tcm_data_outen),       //      .data_outen
		.tcs_tcm_data_in          (generic_tristate_controller_0_tcm_data_in),          //      .data_in
		.tcs_tcm_chipselect_n_out (generic_tristate_controller_0_tcm_chipselect_n_out), //      .chipselect_n_out
		.tcm_address_out          (tristate_conduit_bridge_0_out_tcm_address_out),      //   out.tcm_address_out
		.tcm_read_n_out           (tristate_conduit_bridge_0_out_tcm_read_n_out),       //      .tcm_read_n_out
		.tcm_write_n_out          (tristate_conduit_bridge_0_out_tcm_write_n_out),      //      .tcm_write_n_out
		.tcm_data_out             (tristate_conduit_bridge_0_out_tcm_data_out),         //      .tcm_data_out
		.tcm_chipselect_n_out     (tristate_conduit_bridge_0_out_tcm_chipselect_n_out)  //      .tcm_chipselect_n_out
	);

	nios_system_video_alpha_blender_0 video_alpha_blender_0 (
		.clk                      (clk_clk),                                                            //                    clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                  reset.reset
		.foreground_data          (video_character_buffer_with_dma_0_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),         //                       .ready
		.background_data          (video_rgb_resampler_0_avalon_rgb_source_data),                       // avalon_background_sink.data
		.background_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),              //                       .startofpacket
		.background_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),                //                       .endofpacket
		.background_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),                      //                       .valid
		.background_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),                      //                       .ready
		.output_ready             (video_alpha_blender_0_avalon_blended_source_ready),                  //  avalon_blended_source.ready
		.output_data              (video_alpha_blender_0_avalon_blended_source_data),                   //                       .data
		.output_startofpacket     (video_alpha_blender_0_avalon_blended_source_startofpacket),          //                       .startofpacket
		.output_endofpacket       (video_alpha_blender_0_avalon_blended_source_endofpacket),            //                       .endofpacket
		.output_valid             (video_alpha_blender_0_avalon_blended_source_valid)                   //                       .valid
	);

	nios_system_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (clk_clk),                                                                                  //                       clk.clk
		.reset                (rst_controller_reset_out_reset),                                                           //                     reset.reset
		.ctrl_address         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                 //                          .data
	);

	nios_system_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (clk_clk),                                                         //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                                  //         reset_stream_in.reset
		.clk_stream_out           (clk_0_clk),                                                       //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (video_alpha_blender_0_avalon_blended_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_alpha_blender_0_avalon_blended_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (video_alpha_blender_0_avalon_blended_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (video_alpha_blender_0_avalon_blended_source_valid),               //                        .valid
		.stream_in_data           (video_alpha_blender_0_avalon_blended_source_data),                //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_video_pixel_buffer_dma_0 video_pixel_buffer_dma_0 (
		.clk                  (clk_clk),                                                                    //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                             //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data)                           //                        .data
	);

	nios_system_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                                    //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                             //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_0_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_0_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_0_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)                //                  .data
	);

	nios_system_video_vga_controller_0 video_vga_controller_0 (
		.clk           (clk_0_clk),                                                       //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (video_vga_controller_0_external_interface_CLK),                   // external_interface.export
		.VGA_HS        (video_vga_controller_0_external_interface_HS),                    //                   .export
		.VGA_VS        (video_vga_controller_0_external_interface_VS),                    //                   .export
		.VGA_BLANK     (video_vga_controller_0_external_interface_BLANK),                 //                   .export
		.VGA_SYNC      (video_vga_controller_0_external_interface_SYNC),                  //                   .export
		.VGA_R         (video_vga_controller_0_external_interface_R),                     //                   .export
		.VGA_G         (video_vga_controller_0_external_interface_G),                     //                   .export
		.VGA_B         (video_vga_controller_0_external_interface_B)                      //                   .export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_qsys_0_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_qsys_0_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_qsys_0_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_qsys_0_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_qsys_0_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_qsys_0_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_qsys_0_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_qsys_0_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_qsys_0_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_qsys_0_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_qsys_0_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (nios2_qsys_0_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (nios2_qsys_0_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_done       (),                                                                          //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                      //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                      //    (terminated)
		.ci_slave_multi_result     (),                                                                          //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                               //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                  //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                  //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                                  //    (terminated)
		.multi_ci_master_clk       (),                                                                          //    (terminated)
		.multi_ci_master_reset     (),                                                                          //    (terminated)
		.multi_ci_master_clken     (),                                                                          //    (terminated)
		.multi_ci_master_reset_req (),                                                                          //    (terminated)
		.multi_ci_master_start     (),                                                                          //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                      //    (terminated)
		.multi_ci_master_dataa     (),                                                                          //    (terminated)
		.multi_ci_master_datab     (),                                                                          //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                      //    (terminated)
		.multi_ci_master_n         (),                                                                          //    (terminated)
		.multi_ci_master_readra    (),                                                                          //    (terminated)
		.multi_ci_master_readrb    (),                                                                          //    (terminated)
		.multi_ci_master_writerc   (),                                                                          //    (terminated)
		.multi_ci_master_a         (),                                                                          //    (terminated)
		.multi_ci_master_b         (),                                                                          //    (terminated)
		.multi_ci_master_c         ()                                                                           //    (terminated)
	);

	nios_system_nios2_qsys_0_custom_instruction_master_comb_xconnect nios2_qsys_0_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_estatus),   //           .estatus
		.ci_master1_dataa    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_dataa),     // ci_master1.dataa
		.ci_master1_datab    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_datab),     //           .datab
		.ci_master1_result   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_result),    //           .result
		.ci_master1_n        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_n),         //           .n
		.ci_master1_readra   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_readra),    //           .readra
		.ci_master1_readrb   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_readrb),    //           .readrb
		.ci_master1_writerc  (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_writerc),   //           .writerc
		.ci_master1_a        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_a),         //           .a
		.ci_master1_b        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_b),         //           .b
		.ci_master1_c        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_c),         //           .c
		.ci_master1_ipending (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_ipending),  //           .ipending
		.ci_master1_estatus  (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_0_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                               // (terminated)
		.ci_master_readra    (),                                                                               // (terminated)
		.ci_master_readrb    (),                                                                               // (terminated)
		.ci_master_writerc   (),                                                                               // (terminated)
		.ci_master_a         (),                                                                               // (terminated)
		.ci_master_b         (),                                                                               // (terminated)
		.ci_master_c         (),                                                                               // (terminated)
		.ci_master_ipending  (),                                                                               // (terminated)
		.ci_master_estatus   (),                                                                               // (terminated)
		.ci_master_clk       (),                                                                               // (terminated)
		.ci_master_clken     (),                                                                               // (terminated)
		.ci_master_reset_req (),                                                                               // (terminated)
		.ci_master_reset     (),                                                                               // (terminated)
		.ci_master_start     (),                                                                               // (terminated)
		.ci_master_done      (1'b0),                                                                           // (terminated)
		.ci_slave_clk        (1'b0),                                                                           // (terminated)
		.ci_slave_clken      (1'b0),                                                                           // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                           // (terminated)
		.ci_slave_reset      (1'b0),                                                                           // (terminated)
		.ci_slave_start      (1'b0),                                                                           // (terminated)
		.ci_slave_done       ()                                                                                // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_0_custom_instruction_master_comb_slave_translator1 (
		.ci_slave_dataa      (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master1_estatus),        //          .estatus
		.ci_master_dataa     (nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_qsys_0_custom_instruction_master_comb_slave_translator1_ci_master_result), //          .result
		.ci_master_n         (),                                                                               // (terminated)
		.ci_master_readra    (),                                                                               // (terminated)
		.ci_master_readrb    (),                                                                               // (terminated)
		.ci_master_writerc   (),                                                                               // (terminated)
		.ci_master_a         (),                                                                               // (terminated)
		.ci_master_b         (),                                                                               // (terminated)
		.ci_master_c         (),                                                                               // (terminated)
		.ci_master_ipending  (),                                                                               // (terminated)
		.ci_master_estatus   (),                                                                               // (terminated)
		.ci_master_clk       (),                                                                               // (terminated)
		.ci_master_clken     (),                                                                               // (terminated)
		.ci_master_reset_req (),                                                                               // (terminated)
		.ci_master_reset     (),                                                                               // (terminated)
		.ci_master_start     (),                                                                               // (terminated)
		.ci_master_done      (1'b0),                                                                           // (terminated)
		.ci_slave_clk        (1'b0),                                                                           // (terminated)
		.ci_slave_clken      (1'b0),                                                                           // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                           // (terminated)
		.ci_slave_reset      (1'b0),                                                                           // (terminated)
		.ci_slave_start      (1'b0),                                                                           // (terminated)
		.ci_slave_done       ()                                                                                // (terminated)
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                          (clk_clk),                                                                                  //                                                   clk_0_clk.clk
		.video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                                           //        video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                                       (nios2_qsys_0_data_master_address),                                                         //                                    nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                                   (nios2_qsys_0_data_master_waitrequest),                                                     //                                                            .waitrequest
		.nios2_qsys_0_data_master_byteenable                                    (nios2_qsys_0_data_master_byteenable),                                                      //                                                            .byteenable
		.nios2_qsys_0_data_master_read                                          (nios2_qsys_0_data_master_read),                                                            //                                                            .read
		.nios2_qsys_0_data_master_readdata                                      (nios2_qsys_0_data_master_readdata),                                                        //                                                            .readdata
		.nios2_qsys_0_data_master_readdatavalid                                 (nios2_qsys_0_data_master_readdatavalid),                                                   //                                                            .readdatavalid
		.nios2_qsys_0_data_master_write                                         (nios2_qsys_0_data_master_write),                                                           //                                                            .write
		.nios2_qsys_0_data_master_writedata                                     (nios2_qsys_0_data_master_writedata),                                                       //                                                            .writedata
		.nios2_qsys_0_data_master_debugaccess                                   (nios2_qsys_0_data_master_debugaccess),                                                     //                                                            .debugaccess
		.nios2_qsys_0_instruction_master_address                                (nios2_qsys_0_instruction_master_address),                                                  //                             nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest                            (nios2_qsys_0_instruction_master_waitrequest),                                              //                                                            .waitrequest
		.nios2_qsys_0_instruction_master_read                                   (nios2_qsys_0_instruction_master_read),                                                     //                                                            .read
		.nios2_qsys_0_instruction_master_readdata                               (nios2_qsys_0_instruction_master_readdata),                                                 //                                                            .readdata
		.nios2_qsys_0_instruction_master_readdatavalid                          (nios2_qsys_0_instruction_master_readdatavalid),                                            //                                                            .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_address               (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                                 //            video_pixel_buffer_dma_0_avalon_pixel_dma_master.address
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest           (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),                             //                                                            .waitrequest
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_read                  (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                                    //                                                            .read
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata              (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                                //                                                            .readdata
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid         (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),                           //                                                            .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock                  (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                                    //                                                            .lock
		.generic_tristate_controller_0_uas_address                              (mm_interconnect_0_generic_tristate_controller_0_uas_address),                              //                           generic_tristate_controller_0_uas.address
		.generic_tristate_controller_0_uas_write                                (mm_interconnect_0_generic_tristate_controller_0_uas_write),                                //                                                            .write
		.generic_tristate_controller_0_uas_read                                 (mm_interconnect_0_generic_tristate_controller_0_uas_read),                                 //                                                            .read
		.generic_tristate_controller_0_uas_readdata                             (mm_interconnect_0_generic_tristate_controller_0_uas_readdata),                             //                                                            .readdata
		.generic_tristate_controller_0_uas_writedata                            (mm_interconnect_0_generic_tristate_controller_0_uas_writedata),                            //                                                            .writedata
		.generic_tristate_controller_0_uas_burstcount                           (mm_interconnect_0_generic_tristate_controller_0_uas_burstcount),                           //                                                            .burstcount
		.generic_tristate_controller_0_uas_byteenable                           (mm_interconnect_0_generic_tristate_controller_0_uas_byteenable),                           //                                                            .byteenable
		.generic_tristate_controller_0_uas_readdatavalid                        (mm_interconnect_0_generic_tristate_controller_0_uas_readdatavalid),                        //                                                            .readdatavalid
		.generic_tristate_controller_0_uas_waitrequest                          (mm_interconnect_0_generic_tristate_controller_0_uas_waitrequest),                          //                                                            .waitrequest
		.generic_tristate_controller_0_uas_lock                                 (mm_interconnect_0_generic_tristate_controller_0_uas_lock),                                 //                                                            .lock
		.generic_tristate_controller_0_uas_debugaccess                          (mm_interconnect_0_generic_tristate_controller_0_uas_debugaccess),                          //                                                            .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                                  //                               jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                                    //                                                            .write
		.jtag_uart_0_avalon_jtag_slave_read                                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                                     //                                                            .read
		.jtag_uart_0_avalon_jtag_slave_readdata                                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                                 //                                                            .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                                //                                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                              //                                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                               //                                                            .chipselect
		.new_sdram_controller_0_s1_address                                      (mm_interconnect_0_new_sdram_controller_0_s1_address),                                      //                                   new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                                        (mm_interconnect_0_new_sdram_controller_0_s1_write),                                        //                                                            .write
		.new_sdram_controller_0_s1_read                                         (mm_interconnect_0_new_sdram_controller_0_s1_read),                                         //                                                            .read
		.new_sdram_controller_0_s1_readdata                                     (mm_interconnect_0_new_sdram_controller_0_s1_readdata),                                     //                                                            .readdata
		.new_sdram_controller_0_s1_writedata                                    (mm_interconnect_0_new_sdram_controller_0_s1_writedata),                                    //                                                            .writedata
		.new_sdram_controller_0_s1_byteenable                                   (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),                                   //                                                            .byteenable
		.new_sdram_controller_0_s1_readdatavalid                                (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),                                //                                                            .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                                  (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),                                  //                                                            .waitrequest
		.new_sdram_controller_0_s1_chipselect                                   (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),                                   //                                                            .chipselect
		.nios2_qsys_0_jtag_debug_module_address                                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),                                 //                              nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write                                   (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),                                   //                                                            .write
		.nios2_qsys_0_jtag_debug_module_read                                    (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),                                    //                                                            .read
		.nios2_qsys_0_jtag_debug_module_readdata                                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),                                //                                                            .readdata
		.nios2_qsys_0_jtag_debug_module_writedata                               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),                               //                                                            .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable                              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),                              //                                                            .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest                             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest),                             //                                                            .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess                             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess),                             //                                                            .debugaccess
		.performance_counter_0_control_slave_address                            (mm_interconnect_0_performance_counter_0_control_slave_address),                            //                         performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write                              (mm_interconnect_0_performance_counter_0_control_slave_write),                              //                                                            .write
		.performance_counter_0_control_slave_readdata                           (mm_interconnect_0_performance_counter_0_control_slave_readdata),                           //                                                            .readdata
		.performance_counter_0_control_slave_writedata                          (mm_interconnect_0_performance_counter_0_control_slave_writedata),                          //                                                            .writedata
		.performance_counter_0_control_slave_begintransfer                      (mm_interconnect_0_performance_counter_0_control_slave_begintransfer),                      //                                                            .begintransfer
		.sram_0_avalon_sram_slave_address                                       (mm_interconnect_0_sram_0_avalon_sram_slave_address),                                       //                                    sram_0_avalon_sram_slave.address
		.sram_0_avalon_sram_slave_write                                         (mm_interconnect_0_sram_0_avalon_sram_slave_write),                                         //                                                            .write
		.sram_0_avalon_sram_slave_read                                          (mm_interconnect_0_sram_0_avalon_sram_slave_read),                                          //                                                            .read
		.sram_0_avalon_sram_slave_readdata                                      (mm_interconnect_0_sram_0_avalon_sram_slave_readdata),                                      //                                                            .readdata
		.sram_0_avalon_sram_slave_writedata                                     (mm_interconnect_0_sram_0_avalon_sram_slave_writedata),                                     //                                                            .writedata
		.sram_0_avalon_sram_slave_byteenable                                    (mm_interconnect_0_sram_0_avalon_sram_slave_byteenable),                                    //                                                            .byteenable
		.sram_0_avalon_sram_slave_readdatavalid                                 (mm_interconnect_0_sram_0_avalon_sram_slave_readdatavalid),                                 //                                                            .readdatavalid
		.timer_0_s1_address                                                     (mm_interconnect_0_timer_0_s1_address),                                                     //                                                  timer_0_s1.address
		.timer_0_s1_write                                                       (mm_interconnect_0_timer_0_s1_write),                                                       //                                                            .write
		.timer_0_s1_readdata                                                    (mm_interconnect_0_timer_0_s1_readdata),                                                    //                                                            .readdata
		.timer_0_s1_writedata                                                   (mm_interconnect_0_timer_0_s1_writedata),                                                   //                                                            .writedata
		.timer_0_s1_chipselect                                                  (mm_interconnect_0_timer_0_s1_chipselect),                                                  //                                                            .chipselect
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //  video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                                                            .write
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                                                            .read
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                                                            .readdata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                                                            .writedata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //                                                            .byteenable
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                                                            .waitrequest
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                                                            .chipselect
		.video_character_buffer_with_dma_0_avalon_char_control_slave_address    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // video_character_buffer_with_dma_0_avalon_char_control_slave.address
		.video_character_buffer_with_dma_0_avalon_char_control_slave_write      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                                                            .write
		.video_character_buffer_with_dma_0_avalon_char_control_slave_read       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                                                            .read
		.video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                                                            .readdata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                                                            .writedata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                                                            .byteenable
		.video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                                                            .chipselect
		.video_pixel_buffer_dma_0_avalon_control_slave_address                  (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),                  //               video_pixel_buffer_dma_0_avalon_control_slave.address
		.video_pixel_buffer_dma_0_avalon_control_slave_write                    (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),                    //                                                            .write
		.video_pixel_buffer_dma_0_avalon_control_slave_read                     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),                     //                                                            .read
		.video_pixel_buffer_dma_0_avalon_control_slave_readdata                 (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),                 //                                                            .readdata
		.video_pixel_buffer_dma_0_avalon_control_slave_writedata                (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),                //                                                            .writedata
		.video_pixel_buffer_dma_0_avalon_control_slave_byteenable               (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable)                //                                                            .byteenable
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                           // reset_in1.reset
		.reset_in2      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_0_reset_n),                           // reset_in0.reset
		.reset_in1      (~reset_reset_n),                             // reset_in1.reset
		.reset_in2      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_0_clk),                                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
