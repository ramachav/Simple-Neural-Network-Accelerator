/**
 *	AcceleratorTopMod.sv
 *
 * 	Created	:	26 Nov 2019, 12:44 PM EST
 * 	Author	:	Abhishek Bhaumick
 * 	
 */


module AcceleratorTopMod (
	input 			clk,		// Clock
	input 			clk_en,	// Clock Enable
	input			rst,		// Asynchronous reset active low

	input [ 7:0]	addressIn,
	input [31:0]	dataIn,

	
);

endmodule