/*************************************************************  
*  Floating Point Adder Testbench							 *
*  ECE 69500R SoC Architecture                               *
*  Simple Neural Network Accelerator                         *
*************************************************************/

module fp_adder_tb();

endmodule // fp_adder_tb 

program test (
	input logic clk,
	output logic n_rst,
	output logic [31:0] A,
	output logic [31:0] B,
	input logic [31:0] O
);

initial begin

end
endprogram