/***********************************************************************************  
*  Single Precision Floating Point Multiplier Testbench                            *
*  ECE 69500R SoC Architecture                                                     *
*  Simple Neural Network Accelerator                                               *
***********************************************************************************/

module fp_multiplier_tb();

endmodule // fp_multiplier_tb

program test (
	input logic clk,
	output logic n_rst,
	output logic [31:0] A,
	output logic [31:0] B,
	input logic [31:0] O
);

initial begin

end
endprogram